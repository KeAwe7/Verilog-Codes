`timescale 1ms/1ms

module delays(
	input a,
	input b,
	output out
);

or #5 o1 (out, a, b);

endmodule 